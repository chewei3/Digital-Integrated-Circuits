library verilog;
use verilog.vl_types.all;
entity AS_tb is
end AS_tb;
