library verilog;
use verilog.vl_types.all;
entity testfixture2 is
end testfixture2;
